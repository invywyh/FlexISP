module lambda_arris_v3lua_line43_10(in0, in1, in2, out);
  input [15:0] in0;
  input [15:0] in1;
  input [15:0] in2;
  output [15:0] out;
  
  wire [15:0] cropSpecial0Node_10_pp_0_0_2 = in0;
  wire [15:0] cropSpecial0Node_10_pp_0_0_1 = in1;
  wire [15:0] cropSpecial0Node_10_pp_0_0_0 = in2;
  wire [15:0] c_0_0 = 16'd16383;
  wire [15:0] c_32767_0 = 16'd16383;
  
  wire [15:0] tap_Green_to_Lum_0 = 16'd16383;
  wire [15:0] tap_Blue_to_Lum_0 = 16'd16383;
  wire [15:0] tap_Red_to_Lum_0 = 16'd16383;
  
  wire [15:0] Wxx_8_0 = c_0_0;
  wire [15:0] lambda_arris_v3lua_line43_46_0 = cropSpecial0Node_10_pp_0_0_0;
  wire [15:0] lambda_arris_v3lua_line43_47_0 = lambda_arris_v3lua_line43_46_0;
  wire [15:0] lambda_arris_v3lua_line43_48_0_PP__0__0 = lambda_arris_v3lua_line43_47_0;
  wire [15:0] lambda_arris_v3lua_line43_48_0_PP__0__1 = tap_Red_to_Lum_0;
  wire [15:0] lambda_arris_v3lua_line43_48_0_PP__1__0;
  MULT_pe lambda_arris_v3lua_line43_10_3_0(.clk(),.c(lambda_arris_v3lua_line43_48_0_PP__1__0), .a(lambda_arris_v3lua_line43_48_0_PP__0__0), .b(lambda_arris_v3lua_line43_48_0_PP__0__1));
  wire [15:0] lambda_arris_v3lua_line43_48_0 = lambda_arris_v3lua_line43_48_0_PP__1__0;
  wire [15:0] lambda_arris_v3lua_line43_40_0 = cropSpecial0Node_10_pp_0_0_1;
  wire [15:0] lambda_arris_v3lua_line43_41_0 = lambda_arris_v3lua_line43_40_0;
  wire [15:0] Resp_17_0 = c_32767_0;
  wire [15:0] lambda_arris_v3lua_line43_51_pack_1 = Resp_17_0;
  wire [15:0] lambda_arris_v3lua_line43_42_0_PP__0__0 = lambda_arris_v3lua_line43_41_0;
  wire [15:0] lambda_arris_v3lua_line43_42_0_PP__0__1 = tap_Green_to_Lum_0;
  wire [15:0] lambda_arris_v3lua_line43_42_0_PP__1__0;
  MULT_pe lambda_arris_v3lua_line43_10_8_0(.clk(),.c(lambda_arris_v3lua_line43_42_0_PP__1__0), .a(lambda_arris_v3lua_line43_42_0_PP__0__0), .b(lambda_arris_v3lua_line43_42_0_PP__0__1));
  wire [15:0] lambda_arris_v3lua_line43_42_0 = lambda_arris_v3lua_line43_42_0_PP__1__0;
  wire [15:0] lambda_arris_v3lua_line43_49_pack_1 = lambda_arris_v3lua_line43_42_0;
  wire [15:0] lambda_arris_v3lua_line43_49_pack_0 = lambda_arris_v3lua_line43_48_0;
  wire [15:0] lambda_arris_v3lua_line43_50_pack_1 = Wxx_8_0;
  wire [15:0] lambda_arris_v3lua_line43_43_0 = cropSpecial0Node_10_pp_0_0_2;
  wire [15:0] lambda_arris_v3lua_line43_44_0 = lambda_arris_v3lua_line43_43_0;
  wire [15:0] lambda_arris_v3lua_line43_45_0_PP__0__0 = lambda_arris_v3lua_line43_44_0;
  wire [15:0] lambda_arris_v3lua_line43_45_0_PP__0__1 = tap_Blue_to_Lum_0;
  wire [15:0] lambda_arris_v3lua_line43_45_0_PP__1__0;
  MULT_pe lambda_arris_v3lua_line43_10_14_0(.clk(),.c(lambda_arris_v3lua_line43_45_0_PP__1__0), .a(lambda_arris_v3lua_line43_45_0_PP__0__0), .b(lambda_arris_v3lua_line43_45_0_PP__0__1));
  wire [15:0] lambda_arris_v3lua_line43_45_0 = lambda_arris_v3lua_line43_45_0_PP__1__0;
  wire [15:0] lambda_arris_v3lua_line43_49_pack_2 = lambda_arris_v3lua_line43_45_0;
  wire [15:0] lambda_arris_v3lua_line43_49_0_PP__0__0 = lambda_arris_v3lua_line43_49_pack_2;
  wire [15:0] lambda_arris_v3lua_line43_49_0_PP__0__1 = lambda_arris_v3lua_line43_49_pack_1;
  wire [15:0] lambda_arris_v3lua_line43_49_0_PP__0__2 = lambda_arris_v3lua_line43_49_pack_0;
  wire [15:0] lambda_arris_v3lua_line43_49_0_PP__0__3 = 32'h0;
  wire [15:0] lambda_arris_v3lua_line43_49_0_PP__1__0;
  ALU_pe lambda_arris_v3lua_line43_10_16_0(.clk(),.c(lambda_arris_v3lua_line43_49_0_PP__1__0), .a(lambda_arris_v3lua_line43_49_0_PP__0__0), .b(lambda_arris_v3lua_line43_49_0_PP__0__1));
  wire [15:0] lambda_arris_v3lua_line43_49_0_PP__1__1;
  ALU_pe lambda_arris_v3lua_line43_10_16_1(.clk(),.c(lambda_arris_v3lua_line43_49_0_PP__1__1), .a(lambda_arris_v3lua_line43_49_0_PP__0__2), .b(lambda_arris_v3lua_line43_49_0_PP__0__3));
  wire [15:0] lambda_arris_v3lua_line43_49_0_PP__2__0;
  ALU_pe lambda_arris_v3lua_line43_10_16_2(.clk(),.c(lambda_arris_v3lua_line43_49_0_PP__2__0), .a(lambda_arris_v3lua_line43_49_0_PP__1__0), .b(lambda_arris_v3lua_line43_49_0_PP__1__1));
  wire [15:0] lambda_arris_v3lua_line43_49_0 = lambda_arris_v3lua_line43_49_0_PP__2__0;
  wire [15:0] lambda_arris_v3lua_line43_50_pack_0 = lambda_arris_v3lua_line43_49_0;
  wire [15:0] lambda_arris_v3lua_line43_50_0_PP__0__0 = lambda_arris_v3lua_line43_50_pack_1;
  wire [15:0] lambda_arris_v3lua_line43_50_0_PP__0__1 = lambda_arris_v3lua_line43_50_pack_0;
  wire [15:0] lambda_arris_v3lua_line43_50_0_PP__1__0;
  COMPARE_pe lambda_arris_v3lua_line43_10_18_0(.clk(),.c(lambda_arris_v3lua_line43_50_0_PP__1__0), .a(lambda_arris_v3lua_line43_50_0_PP__0__0), .b(lambda_arris_v3lua_line43_50_0_PP__0__1));
  wire [15:0] lambda_arris_v3lua_line43_50_0 = lambda_arris_v3lua_line43_50_0_PP__1__0;
  wire [15:0] lambda_arris_v3lua_line43_51_pack_0 = lambda_arris_v3lua_line43_50_0;
  wire [15:0] lambda_arris_v3lua_line43_51_0_PP__0__0 = lambda_arris_v3lua_line43_51_pack_1;
  wire [15:0] lambda_arris_v3lua_line43_51_0_PP__0__1 = lambda_arris_v3lua_line43_51_pack_0;
  wire [15:0] lambda_arris_v3lua_line43_51_0_PP__1__0;
  COMPARE_pe lambda_arris_v3lua_line43_10_20_0(.clk(),.c(lambda_arris_v3lua_line43_51_0_PP__1__0), .a(lambda_arris_v3lua_line43_51_0_PP__0__0), .b(lambda_arris_v3lua_line43_51_0_PP__0__1));
  wire [15:0] lambda_arris_v3lua_line43_51_0 = lambda_arris_v3lua_line43_51_0_PP__1__0;
  assign out = lambda_arris_v3lua_line43_51_0;
endmodule // END lambda_arris_v3lua_line43_10


module Resp_5(in0, in1, in2, in3, in4, in5, in6, in7, in8, out);
  input [15:0] in0;
  input [15:0] in1;
  input [15:0] in2;
  input [15:0] in3;
  input [15:0] in4;
  input [15:0] in5;
  input [15:0] in6;
  input [15:0] in7;
  input [15:0] in8;
  output [15:0] out;
  
  wire [15:0] downCast_38_pp_2_2 = in0;
  wire [15:0] downCast_38_pp_2_1 = in1;
  wire [15:0] downCast_38_pp_2_0 = in2;
  wire [15:0] downCast_38_pp_1_2 = in3;
  wire [15:0] downCast_38_pp_1_1 = in4;
  wire [15:0] downCast_38_pp_1_0 = in5;
  wire [15:0] downCast_38_pp_0_2 = in6;
  wire [15:0] downCast_38_pp_0_1 = in7;
  wire [15:0] downCast_38_pp_0_0 = in8;
  wire [15:0] c_1_0 = 16'd16383;
  wire [15:0] c_32767_0 = 16'd16383;
  wire [15:0] c_16_0 = 16'd16383;
  wire [15:0] c_15_0 = 16'd16383;
  
  wire [15:0] tap_K_0 = 16'd16383;
  
  wire [15:0] in1_29_0 = downCast_38_pp_2_0;
  wire [15:0] in1y_22_pack_5 = in1_29_0;
  wire [15:0] in1_31_0 = downCast_38_pp_1_2;
  wire [15:0] in1_26_0 = downCast_38_pp_0_1;
  wire [15:0] in1_27_0 = downCast_38_pp_0_0;
  wire [15:0] in1y_22_pack_3 = in1_27_0;
  wire [15:0] Resp_22_0 = c_32767_0;
  wire [15:0] Wxx_24_pack_1 = Resp_22_0;
  wire [15:0] Resp_31_pack_1 = Resp_22_0;
  wire [15:0] Wyy_19_pack_1 = Resp_22_0;
  wire [15:0] Resp_23_0;
  ALU_pe Resp_5_10_0(.clk(), .c(Resp_23_0), .a(Resp_22_0) ,.b(16'h0));
  wire [15:0] Wxy_15_pack_1 = Resp_23_0;
  wire [15:0] Resp_30_pack_1 = Resp_23_0;
  wire [15:0] in1x_33_0;
  ALU_pe Resp_5_13_0(.clk(), .c(in1x_33_0), .a(in1_27_0) ,.b(16'h0));
  wire [15:0] Wxx_11_0 = c_16_0;
  wire [15:0] in1x_12_0 = c_1_0;
  wire [15:0] in1x_31_0;
  SHIFT_pe Resp_5_16_0(.clk(), .c(in1x_31_0), .a(in1_26_0) ,.b(in1x_12_0));
  wire [15:0] in1_32_0 = downCast_38_pp_1_0;
  wire [15:0] Wxy_16_pack_1 = Resp_22_0;
  wire [15:0] TrSq_9_0 = c_15_0;
  wire [15:0] in1x_36_pack_2 = in1x_33_0;
  wire [15:0] in1_28_0 = downCast_38_pp_2_2;
  wire [15:0] in1x_38_pack_1 = Resp_22_0;
  wire [15:0] in1x_37_pack_1 = Resp_23_0;
  wire [15:0] in1_30_0 = downCast_38_pp_2_1;
  wire [15:0] in1x_35_0;
  SHIFT_pe Resp_5_25_0(.clk(), .c(in1x_35_0), .a(in1_30_0) ,.b(in1x_12_0));
  wire [15:0] in1x_36_pack_4 = in1x_35_0;
  wire [15:0] in1x_36_pack_5 = in1_29_0;
  wire [15:0] in1y_23_pack_1 = Resp_23_0;
  wire [15:0] in1x_32_0;
  ALU_pe Resp_5_29_0(.clk(), .c(in1x_32_0), .a(in1x_31_0) ,.b(16'h0));
  wire [15:0] in1x_36_pack_1 = in1x_32_0;
  wire [15:0] in1y_21_0;
  SHIFT_pe Resp_5_31_0(.clk(), .c(in1y_21_0), .a(in1_32_0) ,.b(in1x_12_0));
  wire [15:0] in1y_22_pack_4 = in1y_21_0;
  wire [15:0] in1x_36_pack_3 = in1_28_0;
  wire [15:0] in1_25_0 = downCast_38_pp_0_2;
  wire [15:0] in1y_19_0;
  SHIFT_pe Resp_5_35_0(.clk(), .c(in1y_19_0), .a(in1_31_0) ,.b(in1x_12_0));
  wire [15:0] in1y_24_pack_1 = Resp_22_0;
  wire [15:0] in1x_30_0;
  ALU_pe Resp_5_37_0(.clk(), .c(in1x_30_0), .a(in1_25_0) ,.b(16'h0));
  wire [15:0] in1x_36_pack_0 = in1x_30_0;
  wire [15:0] in1x_36_0_PP__0__0 = in1x_36_pack_5;
  wire [15:0] in1x_36_0_PP__0__1 = in1x_36_pack_4;
  wire [15:0] in1x_36_0_PP__0__2 = in1x_36_pack_3;
  wire [15:0] in1x_36_0_PP__0__3 = in1x_36_pack_2;
  wire [15:0] in1x_36_0_PP__0__4 = in1x_36_pack_1;
  wire [15:0] in1x_36_0_PP__0__5 = in1x_36_pack_0;
  wire [15:0] in1x_36_0_PP__1__0;
  ALU_pe Resp_5_39_0(.clk(),.c(in1x_36_0_PP__1__0), .a(in1x_36_0_PP__0__0), .b(in1x_36_0_PP__0__1));
  wire [15:0] in1x_36_0_PP__1__1;
  ALU_pe Resp_5_39_1(.clk(),.c(in1x_36_0_PP__1__1), .a(in1x_36_0_PP__0__2), .b(in1x_36_0_PP__0__3));
  wire [15:0] in1x_36_0_PP__1__2;
  ALU_pe Resp_5_39_2(.clk(),.c(in1x_36_0_PP__1__2), .a(in1x_36_0_PP__0__4), .b(in1x_36_0_PP__0__5));
  wire [15:0] in1x_36_0_PP__1__3 = 32'h0;
  wire [15:0] in1x_36_0_PP__2__0;
  ALU_pe Resp_5_39_3(.clk(),.c(in1x_36_0_PP__2__0), .a(in1x_36_0_PP__1__0), .b(in1x_36_0_PP__1__1));
  wire [15:0] in1x_36_0_PP__2__1;
  ALU_pe Resp_5_39_4(.clk(),.c(in1x_36_0_PP__2__1), .a(in1x_36_0_PP__1__2), .b(in1x_36_0_PP__1__3));
  wire [15:0] in1x_36_0_PP__3__0;
  ALU_pe Resp_5_39_5(.clk(),.c(in1x_36_0_PP__3__0), .a(in1x_36_0_PP__2__0), .b(in1x_36_0_PP__2__1));
  wire [15:0] in1x_36_0 = in1x_36_0_PP__3__0;
  wire [15:0] in1x_37_pack_0 = in1x_36_0;
  wire [15:0] in1y_22_pack_0 = in1x_30_0;
  wire [15:0] in1x_34_0;
  ALU_pe Resp_5_42_0(.clk(), .c(in1x_34_0), .a(in1_28_0) ,.b(16'h0));
  wire [15:0] in1y_22_pack_2 = in1x_34_0;
  wire [15:0] Wxx_23_pack_1 = Resp_23_0;
  wire [15:0] Wyy_18_pack_1 = Resp_23_0;
  wire [15:0] in1x_37_0_PP__0__0 = in1x_37_pack_1;
  wire [15:0] in1x_37_0_PP__0__1 = in1x_37_pack_0;
  wire [15:0] in1x_37_0_PP__1__0;
  COMPARE_pe Resp_5_46_0(.clk(),.c(in1x_37_0_PP__1__0), .a(in1x_37_0_PP__0__0), .b(in1x_37_0_PP__0__1));
  wire [15:0] in1x_37_0 = in1x_37_0_PP__1__0;
  wire [15:0] in1x_38_pack_0 = in1x_37_0;
  wire [15:0] in1x_38_0_PP__0__0 = in1x_38_pack_1;
  wire [15:0] in1x_38_0_PP__0__1 = in1x_38_pack_0;
  wire [15:0] in1x_38_0_PP__1__0;
  COMPARE_pe Resp_5_48_0(.clk(),.c(in1x_38_0_PP__1__0), .a(in1x_38_0_PP__0__0), .b(in1x_38_0_PP__0__1));
  wire [15:0] in1x_38_0 = in1x_38_0_PP__1__0;
  wire [15:0] sobel_3_0 = in1x_38_0;
  wire [15:0] Wxx_20_0 = sobel_3_0;
  wire [15:0] Wxx_21_0_PP__0__0 = Wxx_20_0;
  wire [15:0] Wxx_21_0_PP__0__1 = Wxx_20_0;
  wire [15:0] Wxx_21_0_PP__1__0;
  MULT_pe Resp_5_51_0(.clk(),.c(Wxx_21_0_PP__1__0), .a(Wxx_21_0_PP__0__0), .b(Wxx_21_0_PP__0__1));
  wire [15:0] Wxx_21_0 = Wxx_21_0_PP__1__0;
  wire [15:0] Wxx_22_0;
  SHIFT_pe Resp_5_52_0(.clk(), .c(Wxx_22_0), .a(Wxx_21_0) ,.b(Wxx_11_0));
  wire [15:0] Wxx_23_pack_0 = Wxx_22_0;
  wire [15:0] Wxx_23_0_PP__0__0 = Wxx_23_pack_1;
  wire [15:0] Wxx_23_0_PP__0__1 = Wxx_23_pack_0;
  wire [15:0] Wxx_23_0_PP__1__0;
  COMPARE_pe Resp_5_54_0(.clk(),.c(Wxx_23_0_PP__1__0), .a(Wxx_23_0_PP__0__0), .b(Wxx_23_0_PP__0__1));
  wire [15:0] Wxx_23_0 = Wxx_23_0_PP__1__0;
  wire [15:0] Wxx_24_pack_0 = Wxx_23_0;
  wire [15:0] Wxx_24_0_PP__0__0 = Wxx_24_pack_1;
  wire [15:0] Wxx_24_0_PP__0__1 = Wxx_24_pack_0;
  wire [15:0] Wxx_24_0_PP__1__0;
  COMPARE_pe Resp_5_56_0(.clk(),.c(Wxx_24_0_PP__1__0), .a(Wxx_24_0_PP__0__0), .b(Wxx_24_0_PP__0__1));
  wire [15:0] Wxx_24_0 = Wxx_24_0_PP__1__0;
  wire [15:0] in1y_20_0;
  ALU_pe Resp_5_57_0(.clk(), .c(in1y_20_0), .a(in1y_19_0) ,.b(16'h0));
  wire [15:0] in1y_22_pack_1 = in1y_20_0;
  wire [15:0] in1y_22_0_PP__0__0 = in1y_22_pack_5;
  wire [15:0] in1y_22_0_PP__0__1 = in1y_22_pack_4;
  wire [15:0] in1y_22_0_PP__0__2 = in1y_22_pack_3;
  wire [15:0] in1y_22_0_PP__0__3 = in1y_22_pack_2;
  wire [15:0] in1y_22_0_PP__0__4 = in1y_22_pack_1;
  wire [15:0] in1y_22_0_PP__0__5 = in1y_22_pack_0;
  wire [15:0] in1y_22_0_PP__1__0;
  ALU_pe Resp_5_59_0(.clk(),.c(in1y_22_0_PP__1__0), .a(in1y_22_0_PP__0__0), .b(in1y_22_0_PP__0__1));
  wire [15:0] in1y_22_0_PP__1__1;
  ALU_pe Resp_5_59_1(.clk(),.c(in1y_22_0_PP__1__1), .a(in1y_22_0_PP__0__2), .b(in1y_22_0_PP__0__3));
  wire [15:0] in1y_22_0_PP__1__2;
  ALU_pe Resp_5_59_2(.clk(),.c(in1y_22_0_PP__1__2), .a(in1y_22_0_PP__0__4), .b(in1y_22_0_PP__0__5));
  wire [15:0] in1y_22_0_PP__1__3 = 32'h0;
  wire [15:0] in1y_22_0_PP__2__0;
  ALU_pe Resp_5_59_3(.clk(),.c(in1y_22_0_PP__2__0), .a(in1y_22_0_PP__1__0), .b(in1y_22_0_PP__1__1));
  wire [15:0] in1y_22_0_PP__2__1;
  ALU_pe Resp_5_59_4(.clk(),.c(in1y_22_0_PP__2__1), .a(in1y_22_0_PP__1__2), .b(in1y_22_0_PP__1__3));
  wire [15:0] in1y_22_0_PP__3__0;
  ALU_pe Resp_5_59_5(.clk(),.c(in1y_22_0_PP__3__0), .a(in1y_22_0_PP__2__0), .b(in1y_22_0_PP__2__1));
  wire [15:0] in1y_22_0 = in1y_22_0_PP__3__0;
  wire [15:0] in1y_23_pack_0 = in1y_22_0;
  wire [15:0] in1y_23_0_PP__0__0 = in1y_23_pack_1;
  wire [15:0] in1y_23_0_PP__0__1 = in1y_23_pack_0;
  wire [15:0] in1y_23_0_PP__1__0;
  COMPARE_pe Resp_5_61_0(.clk(),.c(in1y_23_0_PP__1__0), .a(in1y_23_0_PP__0__0), .b(in1y_23_0_PP__0__1));
  wire [15:0] in1y_23_0 = in1y_23_0_PP__1__0;
  wire [15:0] in1y_24_pack_0 = in1y_23_0;
  wire [15:0] in1y_24_0_PP__0__0 = in1y_24_pack_1;
  wire [15:0] in1y_24_0_PP__0__1 = in1y_24_pack_0;
  wire [15:0] in1y_24_0_PP__1__0;
  COMPARE_pe Resp_5_63_0(.clk(),.c(in1y_24_0_PP__1__0), .a(in1y_24_0_PP__0__0), .b(in1y_24_0_PP__0__1));
  wire [15:0] in1y_24_0 = in1y_24_0_PP__1__0;
  wire [15:0] sobel_3_1 = in1y_24_0;
  wire [15:0] Wyy_15_0 = sobel_3_1;
  wire [15:0] Wxy_13_0_PP__0__0 = Wxx_20_0;
  wire [15:0] Wxy_13_0_PP__0__1 = Wyy_15_0;
  wire [15:0] Wxy_13_0_PP__1__0;
  MULT_pe Resp_5_66_0(.clk(),.c(Wxy_13_0_PP__1__0), .a(Wxy_13_0_PP__0__0), .b(Wxy_13_0_PP__0__1));
  wire [15:0] Wxy_13_0 = Wxy_13_0_PP__1__0;
  wire [15:0] Wyy_16_0_PP__0__0 = Wyy_15_0;
  wire [15:0] Wyy_16_0_PP__0__1 = Wyy_15_0;
  wire [15:0] Wyy_16_0_PP__1__0;
  MULT_pe Resp_5_67_0(.clk(),.c(Wyy_16_0_PP__1__0), .a(Wyy_16_0_PP__0__0), .b(Wyy_16_0_PP__0__1));
  wire [15:0] Wyy_16_0 = Wyy_16_0_PP__1__0;
  wire [15:0] Wxy_14_0;
  SHIFT_pe Resp_5_68_0(.clk(), .c(Wxy_14_0), .a(Wxy_13_0) ,.b(Wxx_11_0));
  wire [15:0] Wxy_15_pack_0 = Wxy_14_0;
  wire [15:0] Wxy_15_0_PP__0__0 = Wxy_15_pack_1;
  wire [15:0] Wxy_15_0_PP__0__1 = Wxy_15_pack_0;
  wire [15:0] Wxy_15_0_PP__1__0;
  COMPARE_pe Resp_5_70_0(.clk(),.c(Wxy_15_0_PP__1__0), .a(Wxy_15_0_PP__0__0), .b(Wxy_15_0_PP__0__1));
  wire [15:0] Wxy_15_0 = Wxy_15_0_PP__1__0;
  wire [15:0] Wxy_16_pack_0 = Wxy_15_0;
  wire [15:0] Wxy_16_0_PP__0__0 = Wxy_16_pack_1;
  wire [15:0] Wxy_16_0_PP__0__1 = Wxy_16_pack_0;
  wire [15:0] Wxy_16_0_PP__1__0;
  COMPARE_pe Resp_5_72_0(.clk(),.c(Wxy_16_0_PP__1__0), .a(Wxy_16_0_PP__0__0), .b(Wxy_16_0_PP__0__1));
  wire [15:0] Wxy_16_0 = Wxy_16_0_PP__1__0;
  wire [15:0] Det_18_0_PP__0__0 = Wxy_16_0;
  wire [15:0] Det_18_0_PP__0__1 = Wxy_16_0;
  wire [15:0] Det_18_0_PP__1__0;
  MULT_pe Resp_5_73_0(.clk(),.c(Det_18_0_PP__1__0), .a(Det_18_0_PP__0__0), .b(Det_18_0_PP__0__1));
  wire [15:0] Det_18_0 = Det_18_0_PP__1__0;
  wire [15:0] Det_19_0;
  SHIFT_pe Resp_5_74_0(.clk(), .c(Det_19_0), .a(Det_18_0) ,.b(in1x_12_0));
  wire [15:0] Wyy_17_0;
  SHIFT_pe Resp_5_75_0(.clk(), .c(Wyy_17_0), .a(Wyy_16_0) ,.b(Wxx_11_0));
  wire [15:0] Wyy_18_pack_0 = Wyy_17_0;
  wire [15:0] Wyy_18_0_PP__0__0 = Wyy_18_pack_1;
  wire [15:0] Wyy_18_0_PP__0__1 = Wyy_18_pack_0;
  wire [15:0] Wyy_18_0_PP__1__0;
  COMPARE_pe Resp_5_77_0(.clk(),.c(Wyy_18_0_PP__1__0), .a(Wyy_18_0_PP__0__0), .b(Wyy_18_0_PP__0__1));
  wire [15:0] Wyy_18_0 = Wyy_18_0_PP__1__0;
  wire [15:0] Wyy_19_pack_0 = Wyy_18_0;
  wire [15:0] Wyy_19_0_PP__0__0 = Wyy_19_pack_1;
  wire [15:0] Wyy_19_0_PP__0__1 = Wyy_19_pack_0;
  wire [15:0] Wyy_19_0_PP__1__0;
  COMPARE_pe Resp_5_79_0(.clk(),.c(Wyy_19_0_PP__1__0), .a(Wyy_19_0_PP__0__0), .b(Wyy_19_0_PP__0__1));
  wire [15:0] Wyy_19_0 = Wyy_19_0_PP__1__0;
  wire [15:0] Det_16_0_PP__0__0 = Wxx_24_0;
  wire [15:0] Det_16_0_PP__0__1 = Wyy_19_0;
  wire [15:0] Det_16_0_PP__1__0;
  MULT_pe Resp_5_80_0(.clk(),.c(Det_16_0_PP__1__0), .a(Det_16_0_PP__0__0), .b(Det_16_0_PP__0__1));
  wire [15:0] Det_16_0 = Det_16_0_PP__1__0;
  wire [15:0] Det_17_0;
  SHIFT_pe Resp_5_81_0(.clk(), .c(Det_17_0), .a(Det_16_0) ,.b(in1x_12_0));
  wire [15:0] TrSq_15_0_PP__0__0 = Wxx_24_0;
  wire [15:0] TrSq_15_0_PP__0__1 = Wyy_19_0;
  wire [15:0] TrSq_15_0_PP__1__0;
  ALU_pe Resp_5_82_0(.clk(),.c(TrSq_15_0_PP__1__0), .a(TrSq_15_0_PP__0__0), .b(TrSq_15_0_PP__0__1));
  wire [15:0] TrSq_15_0 = TrSq_15_0_PP__1__0;
  wire [15:0] TrSq_16_0;
  SHIFT_pe Resp_5_83_0(.clk(), .c(TrSq_16_0), .a(TrSq_15_0) ,.b(in1x_12_0));
  wire [15:0] TrSq_17_0_PP__0__0 = TrSq_16_0;
  wire [15:0] TrSq_17_0_PP__0__1 = TrSq_16_0;
  wire [15:0] TrSq_17_0_PP__1__0;
  MULT_pe Resp_5_84_0(.clk(),.c(TrSq_17_0_PP__1__0), .a(TrSq_17_0_PP__0__0), .b(TrSq_17_0_PP__0__1));
  wire [15:0] TrSq_17_0 = TrSq_17_0_PP__1__0;
  wire [15:0] TrSq_18_0;
  SHIFT_pe Resp_5_85_0(.clk(), .c(TrSq_18_0), .a(TrSq_17_0) ,.b(TrSq_9_0));
  wire [15:0] Resp1_7_0_PP__0__0 = tap_K_0;
  wire [15:0] Resp1_7_0_PP__0__1 = TrSq_18_0;
  wire [15:0] Resp1_7_0_PP__1__0;
  MULT_pe Resp_5_86_0(.clk(),.c(Resp1_7_0_PP__1__0), .a(Resp1_7_0_PP__0__0), .b(Resp1_7_0_PP__0__1));
  wire [15:0] Resp1_7_0 = Resp1_7_0_PP__1__0;
  wire [15:0] Det_20_0_PP__0__0 = Det_17_0;
  wire [15:0] Det_20_0_PP__0__1 = Det_19_0;
  wire [15:0] Det_20_0_PP__1__0;
  ALU_pe Resp_5_87_0(.clk(),.c(Det_20_0_PP__1__0), .a(Det_20_0_PP__0__0), .b(Det_20_0_PP__0__1));
  wire [15:0] Det_20_0 = Det_20_0_PP__1__0;
  wire [15:0] Resp1_8_0_PP__0__0 = Det_20_0;
  wire [15:0] Resp1_8_0_PP__0__1 = Resp1_7_0;
  wire [15:0] Resp1_8_0_PP__1__0;
  ALU_pe Resp_5_88_0(.clk(),.c(Resp1_8_0_PP__1__0), .a(Resp1_8_0_PP__0__0), .b(Resp1_8_0_PP__0__1));
  wire [15:0] Resp1_8_0 = Resp1_8_0_PP__1__0;
  wire [15:0] Resp_30_pack_0 = Resp1_8_0;
  wire [15:0] Resp_30_0_PP__0__0 = Resp_30_pack_1;
  wire [15:0] Resp_30_0_PP__0__1 = Resp_30_pack_0;
  wire [15:0] Resp_30_0_PP__1__0;
  COMPARE_pe Resp_5_90_0(.clk(),.c(Resp_30_0_PP__1__0), .a(Resp_30_0_PP__0__0), .b(Resp_30_0_PP__0__1));
  wire [15:0] Resp_30_0 = Resp_30_0_PP__1__0;
  wire [15:0] Resp_31_pack_0 = Resp_30_0;
  wire [15:0] Resp_31_0_PP__0__0 = Resp_31_pack_1;
  wire [15:0] Resp_31_0_PP__0__1 = Resp_31_pack_0;
  wire [15:0] Resp_31_0_PP__1__0;
  COMPARE_pe Resp_5_92_0(.clk(),.c(Resp_31_0_PP__1__0), .a(Resp_31_0_PP__0__0), .b(Resp_31_0_PP__0__1));
  wire [15:0] Resp_31_0 = Resp_31_0_PP__1__0;
  wire [15:0] Resp_32_0 = Resp_31_0;
  assign out = Resp_32_0;
endmodule // END Resp_5


module scheduledIRNode_28(in0, in1, in2, out);
  input [15:0] in0;
  input [15:0] in1;
  input [15:0] in2;
  output [15:0] out;
  
  wire [15:0] special0_pp_0_0_2 = in0;
  wire [15:0] special0_pp_0_0_1 = in1;
  wire [15:0] special0_pp_0_0_0 = in2;
  
  
  wire [15:0] cropSpecial0Node_10_0 = special0_pp_0_0_0;
  wire [15:0] cropSpecial0Node_10_1 = special0_pp_0_0_1;
  wire [15:0] cropSpecial0Node_10_2 = special0_pp_0_0_2;
  assign out = cropSpecial0Node_10_2;
  assign out = cropSpecial0Node_10_1;
  assign out = cropSpecial0Node_10_0;
endmodule // END scheduledIRNode_28


module downCast_15(in0, in1, in2, in3, in4, out);
  input [15:0] in0;
  input [15:0] in1;
  input [15:0] in2;
  input [15:0] in3;
  input [15:0] in4;
  output [15:0] out;
  
  wire [15:0] downCast_20_pp_4_0 = in0;
  wire [15:0] downCast_20_pp_3_0 = in1;
  wire [15:0] downCast_20_pp_2_0 = in2;
  wire [15:0] downCast_20_pp_1_0 = in3;
  wire [15:0] downCast_20_pp_0_0 = in4;
  wire [15:0] c_32767_0 = 16'd16383;
  
  wire [15:0] tap_G1_0 = 16'd16383;
  wire [15:0] tap_G0_0 = 16'd16383;
  wire [15:0] tap_G2_0 = 16'd16383;
  wire [15:0] tap_G4_0 = 16'd16383;
  wire [15:0] tap_G3_0 = 16'd16383;
  wire [15:0] tap_R_0 = 16'd16383;
  
  wire [15:0] convolve_1_5__68_0 = tap_G2_0;
  wire [15:0] convolve_1_5__72_0 = tap_G3_0;
  wire [15:0] upCast_37_0 = downCast_20_pp_2_0;
  wire [15:0] convolve_1_5__89_0_PP__0__0 = upCast_37_0;
  wire [15:0] convolve_1_5__89_0_PP__0__1 = convolve_1_5__68_0;
  wire [15:0] convolve_1_5__89_0_PP__1__0;
  MULT_pe downCast_15_3_0(.clk(),.c(convolve_1_5__89_0_PP__1__0), .a(convolve_1_5__89_0_PP__0__0), .b(convolve_1_5__89_0_PP__0__1));
  wire [15:0] convolve_1_5__89_0 = convolve_1_5__89_0_PP__1__0;
  wire [15:0] Resp_20_0 = c_32767_0;
  wire [15:0] convolve_1_5__64_0 = tap_G1_0;
  wire [15:0] upCast_39_0 = downCast_20_pp_3_0;
  wire [15:0] convolve_1_5__70_0 = tap_G4_0;
  wire [15:0] convolve_1_5__93_pack_2 = convolve_1_5__89_0;
  wire [15:0] convolve_1_5__75_0 = tap_R_0;
  wire [15:0] Resp_21_0;
  ALU_pe downCast_15_10_0(.clk(), .c(Resp_21_0), .a(Resp_20_0) ,.b(16'h0));
  wire [15:0] upCast_38_0 = downCast_20_pp_4_0;
  wire [15:0] convolve_1_5__90_0_PP__0__0 = upCast_38_0;
  wire [15:0] convolve_1_5__90_0_PP__0__1 = convolve_1_5__70_0;
  wire [15:0] convolve_1_5__90_0_PP__1__0;
  MULT_pe downCast_15_12_0(.clk(),.c(convolve_1_5__90_0_PP__1__0), .a(convolve_1_5__90_0_PP__0__0), .b(convolve_1_5__90_0_PP__0__1));
  wire [15:0] convolve_1_5__90_0 = convolve_1_5__90_0_PP__1__0;
  wire [15:0] convolve_1_5__93_pack_4 = convolve_1_5__90_0;
  wire [15:0] upCast_36_0 = downCast_20_pp_1_0;
  wire [15:0] convolve_1_5__96_pack_1 = Resp_20_0;
  wire [15:0] convolve_1_5__95_pack_1 = Resp_21_0;
  wire [15:0] convolve_1_5__91_0_PP__0__0 = upCast_39_0;
  wire [15:0] convolve_1_5__91_0_PP__0__1 = convolve_1_5__72_0;
  wire [15:0] convolve_1_5__91_0_PP__1__0;
  MULT_pe downCast_15_17_0(.clk(),.c(convolve_1_5__91_0_PP__1__0), .a(convolve_1_5__91_0_PP__0__0), .b(convolve_1_5__91_0_PP__0__1));
  wire [15:0] convolve_1_5__91_0 = convolve_1_5__91_0_PP__1__0;
  wire [15:0] convolve_1_5__93_pack_3 = convolve_1_5__91_0;
  wire [15:0] convolve_1_5__88_0_PP__0__0 = upCast_36_0;
  wire [15:0] convolve_1_5__88_0_PP__0__1 = convolve_1_5__64_0;
  wire [15:0] convolve_1_5__88_0_PP__1__0;
  MULT_pe downCast_15_19_0(.clk(),.c(convolve_1_5__88_0_PP__1__0), .a(convolve_1_5__88_0_PP__0__0), .b(convolve_1_5__88_0_PP__0__1));
  wire [15:0] convolve_1_5__88_0 = convolve_1_5__88_0_PP__1__0;
  wire [15:0] convolve_1_5__93_pack_1 = convolve_1_5__88_0;
  wire [15:0] upCast_40_0 = downCast_20_pp_0_0;
  wire [15:0] convolve_1_5__66_0 = tap_G0_0;
  wire [15:0] convolve_1_5__92_0_PP__0__0 = upCast_40_0;
  wire [15:0] convolve_1_5__92_0_PP__0__1 = convolve_1_5__66_0;
  wire [15:0] convolve_1_5__92_0_PP__1__0;
  MULT_pe downCast_15_23_0(.clk(),.c(convolve_1_5__92_0_PP__1__0), .a(convolve_1_5__92_0_PP__0__0), .b(convolve_1_5__92_0_PP__0__1));
  wire [15:0] convolve_1_5__92_0 = convolve_1_5__92_0_PP__1__0;
  wire [15:0] convolve_1_5__93_pack_0 = convolve_1_5__92_0;
  wire [15:0] convolve_1_5__93_0_PP__0__0 = convolve_1_5__93_pack_4;
  wire [15:0] convolve_1_5__93_0_PP__0__1 = convolve_1_5__93_pack_3;
  wire [15:0] convolve_1_5__93_0_PP__0__2 = convolve_1_5__93_pack_2;
  wire [15:0] convolve_1_5__93_0_PP__0__3 = convolve_1_5__93_pack_1;
  wire [15:0] convolve_1_5__93_0_PP__0__4 = convolve_1_5__93_pack_0;
  wire [15:0] convolve_1_5__93_0_PP__0__5 = 32'h0;
  wire [15:0] convolve_1_5__93_0_PP__1__0;
  ALU_pe downCast_15_25_0(.clk(),.c(convolve_1_5__93_0_PP__1__0), .a(convolve_1_5__93_0_PP__0__0), .b(convolve_1_5__93_0_PP__0__1));
  wire [15:0] convolve_1_5__93_0_PP__1__1;
  ALU_pe downCast_15_25_1(.clk(),.c(convolve_1_5__93_0_PP__1__1), .a(convolve_1_5__93_0_PP__0__2), .b(convolve_1_5__93_0_PP__0__3));
  wire [15:0] convolve_1_5__93_0_PP__1__2;
  ALU_pe downCast_15_25_2(.clk(),.c(convolve_1_5__93_0_PP__1__2), .a(convolve_1_5__93_0_PP__0__4), .b(convolve_1_5__93_0_PP__0__5));
  wire [15:0] convolve_1_5__93_0_PP__1__3 = 32'h0;
  wire [15:0] convolve_1_5__93_0_PP__2__0;
  ALU_pe downCast_15_25_3(.clk(),.c(convolve_1_5__93_0_PP__2__0), .a(convolve_1_5__93_0_PP__1__0), .b(convolve_1_5__93_0_PP__1__1));
  wire [15:0] convolve_1_5__93_0_PP__2__1;
  ALU_pe downCast_15_25_4(.clk(),.c(convolve_1_5__93_0_PP__2__1), .a(convolve_1_5__93_0_PP__1__2), .b(convolve_1_5__93_0_PP__1__3));
  wire [15:0] convolve_1_5__93_0_PP__3__0;
  ALU_pe downCast_15_25_5(.clk(),.c(convolve_1_5__93_0_PP__3__0), .a(convolve_1_5__93_0_PP__2__0), .b(convolve_1_5__93_0_PP__2__1));
  wire [15:0] convolve_1_5__93_0 = convolve_1_5__93_0_PP__3__0;
  wire [15:0] convolve_1_5__94_0;
  SHIFT_pe downCast_15_26_0(.clk(), .c(convolve_1_5__94_0), .a(convolve_1_5__93_0) ,.b(convolve_1_5__75_0));
  wire [15:0] convolve_1_5__95_pack_0 = convolve_1_5__94_0;
  wire [15:0] convolve_1_5__95_0_PP__0__0 = convolve_1_5__95_pack_1;
  wire [15:0] convolve_1_5__95_0_PP__0__1 = convolve_1_5__95_pack_0;
  wire [15:0] convolve_1_5__95_0_PP__1__0;
  COMPARE_pe downCast_15_28_0(.clk(),.c(convolve_1_5__95_0_PP__1__0), .a(convolve_1_5__95_0_PP__0__0), .b(convolve_1_5__95_0_PP__0__1));
  wire [15:0] convolve_1_5__95_0 = convolve_1_5__95_0_PP__1__0;
  wire [15:0] convolve_1_5__96_pack_0 = convolve_1_5__95_0;
  wire [15:0] convolve_1_5__96_0_PP__0__0 = convolve_1_5__96_pack_1;
  wire [15:0] convolve_1_5__96_0_PP__0__1 = convolve_1_5__96_pack_0;
  wire [15:0] convolve_1_5__96_0_PP__1__0;
  COMPARE_pe downCast_15_30_0(.clk(),.c(convolve_1_5__96_0_PP__1__0), .a(convolve_1_5__96_0_PP__0__0), .b(convolve_1_5__96_0_PP__0__1));
  wire [15:0] convolve_1_5__96_0 = convolve_1_5__96_0_PP__1__0;
  wire [15:0] downCast_38_0 = convolve_1_5__96_0;
  assign out = downCast_38_0;
endmodule // END downCast_15


module NMS_10(in0, in1, in2, in3, in4, in5, in6, in7, in8, out);
  input [15:0] in0;
  input [15:0] in1;
  input [15:0] in2;
  input [15:0] in3;
  input [15:0] in4;
  input [15:0] in5;
  input [15:0] in6;
  input [15:0] in7;
  input [15:0] in8;
  output [15:0] out;
  
  wire [15:0] Resp_32_pp_2_2 = in0;
  wire [15:0] Resp_32_pp_2_1 = in1;
  wire [15:0] Resp_32_pp_2_0 = in2;
  wire [15:0] Resp_32_pp_1_2 = in3;
  wire [15:0] Resp_32_pp_1_1 = in4;
  wire [15:0] Resp_32_pp_1_0 = in5;
  wire [15:0] Resp_32_pp_0_2 = in6;
  wire [15:0] Resp_32_pp_0_1 = in7;
  wire [15:0] Resp_32_pp_0_0 = in8;
  wire [15:0] c_0_0 = 16'd16383;
  wire [15:0] c_255_0 = 16'd16383;
  
  wire [15:0] tap_Peak_0 = 16'd16383;
  
  wire [15:0] PE_4_0;
  LOGIC_pe NMS_10_0_0(.clk(), .c(PE_4_0), .a(Resp_32_pp_1_1) ,.b(Resp_32_pp_2_1));
  wire [15:0] NMS_5_0 = c_255_0;
  wire [15:0] P_7_0 = Resp_32_pp_1_1;
  wire [15:0] P_8_0;
  LOGIC_pe NMS_10_3_0(.clk(), .c(P_8_0), .a(P_7_0) ,.b(tap_Peak_0));
  wire [15:0] PS_4_0;
  LOGIC_pe NMS_10_4_0(.clk(), .c(PS_4_0), .a(Resp_32_pp_1_1) ,.b(Resp_32_pp_1_0));
  wire [15:0] PW_4_0;
  LOGIC_pe NMS_10_5_0(.clk(), .c(PW_4_0), .a(Resp_32_pp_1_1) ,.b(Resp_32_pp_0_1));
  wire [15:0] Pk_13_0;
  ALU_pe NMS_10_6_0(.clk(), .c(Pk_13_0), .a(P_8_0) ,.b(PW_4_0));
  wire [15:0] Pk_14_0;
  ALU_pe NMS_10_7_0(.clk(), .c(Pk_14_0), .a(Pk_13_0) ,.b(PE_4_0));
  wire [15:0] Pk_15_0;
  ALU_pe NMS_10_8_0(.clk(), .c(Pk_15_0), .a(Pk_14_0) ,.b(PS_4_0));
  wire [15:0] PN_4_0;
  LOGIC_pe NMS_10_9_0(.clk(), .c(PN_4_0), .a(Resp_32_pp_1_1) ,.b(Resp_32_pp_1_2));
  wire [15:0] Pk_16_0;
  ALU_pe NMS_10_10_0(.clk(), .c(Pk_16_0), .a(Pk_15_0) ,.b(PN_4_0));
  wire [15:0] Wxx_25_0 = c_0_0;
  wire [15:0] NMS_10_0;
  MUX_pe NMS_10_12_0(.clk(), .c(NMS_10_0), .s(Pk_16_0), .a(NMS_5_0) ,.b(Wxx_25_0));
  wire [15:0] NMS_11_0 = NMS_10_0;
  assign out = NMS_11_0;
endmodule // END NMS_10


module downCast_13(in0, in1, in2, in3, in4, out);
  input [15:0] in0;
  input [15:0] in1;
  input [15:0] in2;
  input [15:0] in3;
  input [15:0] in4;
  output [15:0] out;
  
  wire [15:0] lambda_arris_v3lua_line43_51_pp_0_4 = in0;
  wire [15:0] lambda_arris_v3lua_line43_51_pp_0_3 = in1;
  wire [15:0] lambda_arris_v3lua_line43_51_pp_0_2 = in2;
  wire [15:0] lambda_arris_v3lua_line43_51_pp_0_1 = in3;
  wire [15:0] lambda_arris_v3lua_line43_51_pp_0_0 = in4;
  wire [15:0] c_32767_0 = 16'd16383;
  
  wire [15:0] tap_G1_0 = 16'd16383;
  wire [15:0] tap_G0_0 = 16'd16383;
  wire [15:0] tap_G2_0 = 16'd16383;
  wire [15:0] tap_G4_0 = 16'd16383;
  wire [15:0] tap_G3_0 = 16'd16383;
  wire [15:0] tap_R_0 = 16'd16383;
  
  wire [15:0] convolve_1_5__35_0 = tap_G2_0;
  wire [15:0] convolve_1_5__37_0 = tap_G3_0;
  wire [15:0] upCast_22_0 = lambda_arris_v3lua_line43_51_pp_0_2;
  wire [15:0] convolve_1_5__56_0_PP__0__0 = upCast_22_0;
  wire [15:0] convolve_1_5__56_0_PP__0__1 = convolve_1_5__35_0;
  wire [15:0] convolve_1_5__56_0_PP__1__0;
  MULT_pe downCast_13_3_0(.clk(),.c(convolve_1_5__56_0_PP__1__0), .a(convolve_1_5__56_0_PP__0__0), .b(convolve_1_5__56_0_PP__0__1));
  wire [15:0] convolve_1_5__56_0 = convolve_1_5__56_0_PP__1__0;
  wire [15:0] Resp_18_0 = c_32767_0;
  wire [15:0] convolve_1_5__31_0 = tap_G1_0;
  wire [15:0] upCast_24_0 = lambda_arris_v3lua_line43_51_pp_0_1;
  wire [15:0] convolve_1_5__39_0 = tap_G4_0;
  wire [15:0] convolve_1_5__60_pack_2 = convolve_1_5__56_0;
  wire [15:0] convolve_1_5__42_0 = tap_R_0;
  wire [15:0] Resp_19_0;
  ALU_pe downCast_13_10_0(.clk(), .c(Resp_19_0), .a(Resp_18_0) ,.b(16'h0));
  wire [15:0] upCast_23_0 = lambda_arris_v3lua_line43_51_pp_0_0;
  wire [15:0] convolve_1_5__57_0_PP__0__0 = upCast_23_0;
  wire [15:0] convolve_1_5__57_0_PP__0__1 = convolve_1_5__39_0;
  wire [15:0] convolve_1_5__57_0_PP__1__0;
  MULT_pe downCast_13_12_0(.clk(),.c(convolve_1_5__57_0_PP__1__0), .a(convolve_1_5__57_0_PP__0__0), .b(convolve_1_5__57_0_PP__0__1));
  wire [15:0] convolve_1_5__57_0 = convolve_1_5__57_0_PP__1__0;
  wire [15:0] convolve_1_5__60_pack_4 = convolve_1_5__57_0;
  wire [15:0] upCast_21_0 = lambda_arris_v3lua_line43_51_pp_0_3;
  wire [15:0] convolve_1_5__63_pack_1 = Resp_18_0;
  wire [15:0] convolve_1_5__62_pack_1 = Resp_19_0;
  wire [15:0] convolve_1_5__58_0_PP__0__0 = upCast_24_0;
  wire [15:0] convolve_1_5__58_0_PP__0__1 = convolve_1_5__37_0;
  wire [15:0] convolve_1_5__58_0_PP__1__0;
  MULT_pe downCast_13_17_0(.clk(),.c(convolve_1_5__58_0_PP__1__0), .a(convolve_1_5__58_0_PP__0__0), .b(convolve_1_5__58_0_PP__0__1));
  wire [15:0] convolve_1_5__58_0 = convolve_1_5__58_0_PP__1__0;
  wire [15:0] convolve_1_5__60_pack_3 = convolve_1_5__58_0;
  wire [15:0] convolve_1_5__55_0_PP__0__0 = upCast_21_0;
  wire [15:0] convolve_1_5__55_0_PP__0__1 = convolve_1_5__31_0;
  wire [15:0] convolve_1_5__55_0_PP__1__0;
  MULT_pe downCast_13_19_0(.clk(),.c(convolve_1_5__55_0_PP__1__0), .a(convolve_1_5__55_0_PP__0__0), .b(convolve_1_5__55_0_PP__0__1));
  wire [15:0] convolve_1_5__55_0 = convolve_1_5__55_0_PP__1__0;
  wire [15:0] convolve_1_5__60_pack_1 = convolve_1_5__55_0;
  wire [15:0] upCast_25_0 = lambda_arris_v3lua_line43_51_pp_0_4;
  wire [15:0] convolve_1_5__33_0 = tap_G0_0;
  wire [15:0] convolve_1_5__59_0_PP__0__0 = upCast_25_0;
  wire [15:0] convolve_1_5__59_0_PP__0__1 = convolve_1_5__33_0;
  wire [15:0] convolve_1_5__59_0_PP__1__0;
  MULT_pe downCast_13_23_0(.clk(),.c(convolve_1_5__59_0_PP__1__0), .a(convolve_1_5__59_0_PP__0__0), .b(convolve_1_5__59_0_PP__0__1));
  wire [15:0] convolve_1_5__59_0 = convolve_1_5__59_0_PP__1__0;
  wire [15:0] convolve_1_5__60_pack_0 = convolve_1_5__59_0;
  wire [15:0] convolve_1_5__60_0_PP__0__0 = convolve_1_5__60_pack_4;
  wire [15:0] convolve_1_5__60_0_PP__0__1 = convolve_1_5__60_pack_3;
  wire [15:0] convolve_1_5__60_0_PP__0__2 = convolve_1_5__60_pack_2;
  wire [15:0] convolve_1_5__60_0_PP__0__3 = convolve_1_5__60_pack_1;
  wire [15:0] convolve_1_5__60_0_PP__0__4 = convolve_1_5__60_pack_0;
  wire [15:0] convolve_1_5__60_0_PP__0__5 = 32'h0;
  wire [15:0] convolve_1_5__60_0_PP__1__0;
  ALU_pe downCast_13_25_0(.clk(),.c(convolve_1_5__60_0_PP__1__0), .a(convolve_1_5__60_0_PP__0__0), .b(convolve_1_5__60_0_PP__0__1));
  wire [15:0] convolve_1_5__60_0_PP__1__1;
  ALU_pe downCast_13_25_1(.clk(),.c(convolve_1_5__60_0_PP__1__1), .a(convolve_1_5__60_0_PP__0__2), .b(convolve_1_5__60_0_PP__0__3));
  wire [15:0] convolve_1_5__60_0_PP__1__2;
  ALU_pe downCast_13_25_2(.clk(),.c(convolve_1_5__60_0_PP__1__2), .a(convolve_1_5__60_0_PP__0__4), .b(convolve_1_5__60_0_PP__0__5));
  wire [15:0] convolve_1_5__60_0_PP__1__3 = 32'h0;
  wire [15:0] convolve_1_5__60_0_PP__2__0;
  ALU_pe downCast_13_25_3(.clk(),.c(convolve_1_5__60_0_PP__2__0), .a(convolve_1_5__60_0_PP__1__0), .b(convolve_1_5__60_0_PP__1__1));
  wire [15:0] convolve_1_5__60_0_PP__2__1;
  ALU_pe downCast_13_25_4(.clk(),.c(convolve_1_5__60_0_PP__2__1), .a(convolve_1_5__60_0_PP__1__2), .b(convolve_1_5__60_0_PP__1__3));
  wire [15:0] convolve_1_5__60_0_PP__3__0;
  ALU_pe downCast_13_25_5(.clk(),.c(convolve_1_5__60_0_PP__3__0), .a(convolve_1_5__60_0_PP__2__0), .b(convolve_1_5__60_0_PP__2__1));
  wire [15:0] convolve_1_5__60_0 = convolve_1_5__60_0_PP__3__0;
  wire [15:0] convolve_1_5__61_0;
  SHIFT_pe downCast_13_26_0(.clk(), .c(convolve_1_5__61_0), .a(convolve_1_5__60_0) ,.b(convolve_1_5__42_0));
  wire [15:0] convolve_1_5__62_pack_0 = convolve_1_5__61_0;
  wire [15:0] convolve_1_5__62_0_PP__0__0 = convolve_1_5__62_pack_1;
  wire [15:0] convolve_1_5__62_0_PP__0__1 = convolve_1_5__62_pack_0;
  wire [15:0] convolve_1_5__62_0_PP__1__0;
  COMPARE_pe downCast_13_28_0(.clk(),.c(convolve_1_5__62_0_PP__1__0), .a(convolve_1_5__62_0_PP__0__0), .b(convolve_1_5__62_0_PP__0__1));
  wire [15:0] convolve_1_5__62_0 = convolve_1_5__62_0_PP__1__0;
  wire [15:0] convolve_1_5__63_pack_0 = convolve_1_5__62_0;
  wire [15:0] convolve_1_5__63_0_PP__0__0 = convolve_1_5__63_pack_1;
  wire [15:0] convolve_1_5__63_0_PP__0__1 = convolve_1_5__63_pack_0;
  wire [15:0] convolve_1_5__63_0_PP__1__0;
  COMPARE_pe downCast_13_30_0(.clk(),.c(convolve_1_5__63_0_PP__1__0), .a(convolve_1_5__63_0_PP__0__0), .b(convolve_1_5__63_0_PP__0__1));
  wire [15:0] convolve_1_5__63_0 = convolve_1_5__63_0_PP__1__0;
  wire [15:0] downCast_20_0 = convolve_1_5__63_0;
  assign out = downCast_20_0;
endmodule // END downCast_13


module LineBuf(clk,in,out);
input clk;
input [15:0] in;
output [15:0] out;
assign out = in;
endmodule

module top(clk, TOP_in0, TOP_out0);
  input clk;
  input [15:0] TOP_in0;
  output [15:0] TOP_out0;
  
  wire [15:0] LB_TOP_in0_out = TOP_in0;
  wire [15:0] cropSpecial0Node_10;
  wire[15:0] LB_cropSpecial0Node_10_out;
  LineBuf LBcropSpecial0Node_10(.clk(clk), .in(cropSpecial0Node_10), .out(LB_cropSpecial0Node_10_out));
  scheduledIRNode_28 scheduledIRNode_28_0(.in0(LB_TOP_in0_out), .in1(LB_TOP_in0_out), .in2(LB_TOP_in0_out), .out(cropSpecial0Node_10));
  wire [15:0] lambda_arris_v3lua_line43_51;
  wire[15:0] LB_lambda_arris_v3lua_line43_51_out;
  LineBuf LBlambda_arris_v3lua_line43_51(.clk(clk), .in(lambda_arris_v3lua_line43_51), .out(LB_lambda_arris_v3lua_line43_51_out));
  lambda_arris_v3lua_line43_10 lambda_arris_v3lua_line43_10_1(.in0(LB_cropSpecial0Node_10_out), .in1(LB_cropSpecial0Node_10_out), .in2(LB_cropSpecial0Node_10_out), .out(lambda_arris_v3lua_line43_51));
  wire [15:0] downCast_20;
  wire[15:0] LB_downCast_20_out;
  LineBuf LBdownCast_20(.clk(clk), .in(downCast_20), .out(LB_downCast_20_out));
  downCast_13 downCast_13_2(.in0(LB_lambda_arris_v3lua_line43_51_out), .in1(LB_lambda_arris_v3lua_line43_51_out), .in2(LB_lambda_arris_v3lua_line43_51_out), .in3(LB_lambda_arris_v3lua_line43_51_out), .in4(LB_lambda_arris_v3lua_line43_51_out), .out(downCast_20));
  wire [15:0] downCast_38;
  wire[15:0] LB_downCast_38_out;
  LineBuf LBdownCast_38(.clk(clk), .in(downCast_38), .out(LB_downCast_38_out));
  downCast_15 downCast_15_3(.in0(LB_downCast_20_out), .in1(LB_downCast_20_out), .in2(LB_downCast_20_out), .in3(LB_downCast_20_out), .in4(LB_downCast_20_out), .out(downCast_38));
  wire [15:0] Resp_32;
  wire[15:0] LB_Resp_32_out;
  LineBuf LBResp_32(.clk(clk), .in(Resp_32), .out(LB_Resp_32_out));
  Resp_5 Resp_5_4(.in0(LB_downCast_38_out), .in1(LB_downCast_38_out), .in2(LB_downCast_38_out), .in3(LB_downCast_38_out), .in4(LB_downCast_38_out), .in5(LB_downCast_38_out), .in6(LB_downCast_38_out), .in7(LB_downCast_38_out), .in8(LB_downCast_38_out), .out(Resp_32));
  wire [15:0] NMS_11;
  wire[15:0] LB_NMS_11_out;
  LineBuf LBNMS_11(.clk(clk), .in(NMS_11), .out(LB_NMS_11_out));
  NMS_10 NMS_10_5(.in0(LB_Resp_32_out), .in1(LB_Resp_32_out), .in2(LB_Resp_32_out), .in3(LB_Resp_32_out), .in4(LB_Resp_32_out), .in5(LB_Resp_32_out), .in6(LB_Resp_32_out), .in7(LB_Resp_32_out), .in8(LB_Resp_32_out), .out(NMS_11));
  assign TOP_out0 = LB_NMS_11_out;
endmodule
